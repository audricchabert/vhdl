 entity regn is
 generic (N : natural :=16 ); 
 port(insn_in);
 end regn;
 
 architecture regna of regn is
 begin
 
 
 
 end regna;